`include "NOR1.v"
module NOR_tb;
  reg a;
  reg b;
  wire c;
  NOR1 uut(.a(a),.b(b),.c(c));
  initial
    begin
      $dumpfile("NOR_tb.vcd");
      $dumpvars(0,NOR_tb);
      a=0;
      b=0;
      #100;
      a=0;
      b=1;
      #100;
      a=1;
      b=0;
      #100;
      a=1;
      b=1;
      #100;
    end
endmodule